`define  ETRACE_CFG       6'd0  //configuration
`define  ETRACE_REGS      4'hF  //group decode
`define  ETRACE_MEM       4'hA  //group decode
