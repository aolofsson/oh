module BUFIO (/*AUTOARG*/
   // Outputs
   O,
   // Inputs
   I
   );

   output O;
   input  I;
    
   assign O=I;
     
endmodule
