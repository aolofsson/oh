module oh_hamming_enc (/*AUTOARG*/
   // Outputs
   out,
   // Inputs
   in, reset
   );

   output out;

   input in;
   input reset;
endmodule // oh_hamming_enc


