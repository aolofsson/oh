`ifndef GPIO_REGMAP_VH_
 `define GPIO_REGMAP_VH_
 `define GPIO_OEN      6'h0
 `define GPIO_OUT      6'h2
 `define GPIO_IEN      6'h4
 `define GPIO_IN       6'h6
 `define GPIO_OUTAND   6'h8
 `define GPIO_OUTORR   6'ha
 `define GPIO_OUTXOR   6'hc
 `define GPIO_IRQMASK  6'he
`endif
