module oh_8b10b_decode (/*AUTOINST*/);

endmodule // oh_pll
