`define CFG_TARGET "GENERIC"
`define CFG_RANDOM "1"
