module BUFIO (/*AUTOARG*/
   // Outputs
   O,
   // Inputs
   I
   );
   input I;
   output O;

   assign O=I;
   
endmodule // BUFIO

