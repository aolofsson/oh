module oh_ecc_read (/*AUTOARG*/);


endmodule // oh_ecc_read

