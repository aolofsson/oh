module oh_hamming_enc (/*AUTOARG*/
   // Outputs
   out,
   // Inputs
   in, reset
   );

 
endmodule // oh_hamming_enc


