//#############################################################################
//# Function: Charge Keeper Cell                                              #
//# Copyright: OH Project Authors. ALl rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_keeper
   (
    inout z
    );

endmodule
