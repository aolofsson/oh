//#############################################################################
//# Function: Decap Cell                                                      #
//# Copyright: OH Project Authors. ALl rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_decap #(parameter PROP = "DEFAULT")   (
    input  vss,
    output vdd
    );

endmodule
