//#############################################################################
//# Function: Isolation buffer for multi supply domains                       #
//#############################################################################
//# Author:   Andreas Olofsson                                                #
//# License:  MIT (see below)                                                 # 
//#############################################################################

module oh_pwr_isolate (/*AUTOARG*/
   // Outputs
   out,
   // Inputs
   vdd, vss, niso, in
   );

   parameter       DW=1;  // width of macro

   input           vdd;    // supply (set to 1 if valid)
   input           vss;    // ground (set to 0 if valid)
   input 	   niso;   // active low isolation signal
   input [DW-1:0]  in;     // input signal
   output [DW-1:0] out;    // buffered output signal
   
`ifdef TARGET_SIM   
   assign out[DW-1:0] = ((vdd===1'b1) && (vss===1'b0)) ? ({(DW){niso}} & in[DW-1:0]):
		                                         {(DW){1'bX}};
`else
   assign out[DW-1:0] = {(DW){niso}} & in[DW-1:0];
`endif
   
endmodule // oh_buf

///////////////////////////////////////////////////////////////////////////////
// The MIT License (MIT)                                                     //
//                                                                           //
// Copyright (c) 2015-2016, Adapteva, Inc.                                   //
//                                                                           //
// Permission is hereby granted, free of charge, to any person obtaining a   //
// copy of this software and associated documentation files (the "Software") //
// to deal in the Software without restriction, including without limitation // 
// the rights to use, copy, modify, merge, publish, distribute, sublicense,  //
// and/or sell copies of the Software, and to permit persons to whom the     //
// Software is furnished to do so, subject to the following conditions:      //
//                                                                           //
// The above copyright notice and this permission notice shall be included   // 
// in all copies or substantial portions of the Software.                    //
//                                                                           //
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS   //
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF                //
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.    //
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY      //
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT //
// OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR  //
// THE USE OR OTHER DEALINGS IN THE SOFTWARE.                                //
//                                                                           // 
///////////////////////////////////////////////////////////////////////////////
