
module OBUFT (O, I, T);

    parameter CAPACITANCE = "DONT_CARE";
    parameter integer DRIVE = 12;
    parameter IOSTANDARD = "DEFAULT";


   output 	      O;
   input 	      I, T;

   
endmodule

