//#############################################################################
//# Function: Antenna Diode                                                   #
//# Copyright: OH Project Authors. ALl rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_antenna #(parameter PROP = "DEFAULT")   (
    input  vss,
    output z
    );

endmodule
