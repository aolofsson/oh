//Version v5_5
module processing_system7 (
  #(
  parameter integer C_USE_DEFAULT_ACP_USER_VAL = 1,
  parameter integer C_S_AXI_ACP_ARUSER_VAL = 31,
  parameter integer C_S_AXI_ACP_AWUSER_VAL = 31,
  parameter integer C_M_AXI_GP0_THREAD_ID_WIDTH = 12,
  parameter integer C_M_AXI_GP1_THREAD_ID_WIDTH = 12, 
  parameter integer C_M_AXI_GP0_ENABLE_STATIC_REMAP = 1,
  parameter integer C_M_AXI_GP1_ENABLE_STATIC_REMAP = 1, 
  parameter integer C_M_AXI_GP0_ID_WIDTH = 12,
  parameter integer C_M_AXI_GP1_ID_WIDTH = 12,
  parameter integer C_S_AXI_GP0_ID_WIDTH = 6,
  parameter integer C_S_AXI_GP1_ID_WIDTH = 6,
  parameter integer C_S_AXI_HP0_ID_WIDTH = 6,
  parameter integer C_S_AXI_HP1_ID_WIDTH = 6,
  parameter integer C_S_AXI_HP2_ID_WIDTH = 6,
  parameter integer C_S_AXI_HP3_ID_WIDTH = 6,
  parameter integer C_S_AXI_ACP_ID_WIDTH = 3,
  parameter integer C_S_AXI_HP0_DATA_WIDTH = 64,
  parameter integer C_S_AXI_HP1_DATA_WIDTH = 64,
  parameter integer C_S_AXI_HP2_DATA_WIDTH = 64,
  parameter integer C_S_AXI_HP3_DATA_WIDTH = 64,
  parameter integer C_INCLUDE_ACP_TRANS_CHECK = 0,
  parameter integer C_NUM_F2P_INTR_INPUTS = 1,
  parameter         C_FCLK_CLK0_BUF = "TRUE",
  parameter         C_FCLK_CLK1_BUF = "TRUE",
  parameter         C_FCLK_CLK2_BUF = "TRUE",
  parameter         C_FCLK_CLK3_BUF = "TRUE",
  parameter integer C_EMIO_GPIO_WIDTH = 64,
  parameter integer C_INCLUDE_TRACE_BUFFER = 0,
  parameter integer C_TRACE_BUFFER_FIFO_SIZE = 128,
  parameter integer C_TRACE_BUFFER_CLOCK_DELAY = 12,
  parameter integer USE_TRACE_DATA_EDGE_DETECTOR = 0,
  parameter integer C_TRACE_PIPELINE_WIDTH = 8,
  parameter         C_PS7_SI_REV = "PRODUCTION",
  parameter integer C_EN_EMIO_ENET0 = 0,
  parameter integer C_EN_EMIO_ENET1 = 0,
  parameter integer C_EN_EMIO_TRACE = 0,
  parameter integer C_DQ_WIDTH = 32,
  parameter integer C_DQS_WIDTH = 4,
  parameter integer C_DM_WIDTH = 4,
  parameter integer C_MIO_PRIMITIVE = 54,
  parameter	    C_PACKAGE_NAME = "clg484",
  parameter         C_IRQ_F2P_MODE = "DIRECT",
  parameter         C_TRACE_INTERNAL_WIDTH = 32,
  parameter integer C_EN_EMIO_PJTAG = 0
) 
  //FMIO CAN0
  output 				       CAN0_PHY_TX,
  input 				       CAN0_PHY_RX,

  //FMIO CAN1
  output 				       CAN1_PHY_TX, 
  input 				       CAN1_PHY_RX,
  
  //FMIO ENET0
  output reg 				       ENET0_GMII_TX_EN,
  output reg 				       ENET0_GMII_TX_ER,
  output 				       ENET0_MDIO_MDC,
  output 				       ENET0_MDIO_O,
  output 				       ENET0_MDIO_T,
  output 				       ENET0_PTP_DELAY_REQ_RX,
  output 				       ENET0_PTP_DELAY_REQ_TX,
  output 				       ENET0_PTP_PDELAY_REQ_RX,
  output 				       ENET0_PTP_PDELAY_REQ_TX,
  output 				       ENET0_PTP_PDELAY_RESP_RX,
  output 				       ENET0_PTP_PDELAY_RESP_TX,
  output 				       ENET0_PTP_SYNC_FRAME_RX,
  output 				       ENET0_PTP_SYNC_FRAME_TX,
  output 				       ENET0_SOF_RX,
  output 				       ENET0_SOF_TX,
  
  
  output reg [7:0] 			       ENET0_GMII_TXD, 

  
  input 				       ENET0_GMII_COL,
  input 				       ENET0_GMII_CRS,
  input 				       ENET0_GMII_RX_CLK,
  input 				       ENET0_GMII_RX_DV,
  input 				       ENET0_GMII_RX_ER,
  input 				       ENET0_GMII_TX_CLK,
  input 				       ENET0_MDIO_I,
  input 				       ENET0_EXT_INTIN,
  input [7:0] 				       ENET0_GMII_RXD, 

  //FMIO ENET1
  output reg 				       ENET1_GMII_TX_EN,
  output reg 				       ENET1_GMII_TX_ER,
  output 				       ENET1_MDIO_MDC,
  output 				       ENET1_MDIO_O,
  output 				       ENET1_MDIO_T,
  output 				       ENET1_PTP_DELAY_REQ_RX,
  output 				       ENET1_PTP_DELAY_REQ_TX,
  output 				       ENET1_PTP_PDELAY_REQ_RX,
  output 				       ENET1_PTP_PDELAY_REQ_TX,
  output 				       ENET1_PTP_PDELAY_RESP_RX,
  output 				       ENET1_PTP_PDELAY_RESP_TX,
  output 				       ENET1_PTP_SYNC_FRAME_RX,
  output 				       ENET1_PTP_SYNC_FRAME_TX,
  output 				       ENET1_SOF_RX,
  output 				       ENET1_SOF_TX,
  output reg [7:0] 			       ENET1_GMII_TXD, 

  input 				       ENET1_GMII_COL,
  input 				       ENET1_GMII_CRS,
  input 				       ENET1_GMII_RX_CLK,
  input 				       ENET1_GMII_RX_DV,
  input 				       ENET1_GMII_RX_ER,
  input 				       ENET1_GMII_TX_CLK,
  input 				       ENET1_MDIO_I,
  input 				       ENET1_EXT_INTIN, 
  input [7:0] 				       ENET1_GMII_RXD,
  
  //FMIO GPIO
  input [(C_EMIO_GPIO_WIDTH-1):0] 	       GPIO_I,
  output [(C_EMIO_GPIO_WIDTH-1):0] 	       GPIO_O,
  output [(C_EMIO_GPIO_WIDTH-1):0] 	       GPIO_T, 
  
  //FMIO I2C0
  input 				       I2C0_SDA_I,
  output 				       I2C0_SDA_O,
  output 				       I2C0_SDA_T,
  input 				       I2C0_SCL_I,
  output 				       I2C0_SCL_O,
  output 				       I2C0_SCL_T,

  //FMIO I2C1
  input 				       I2C1_SDA_I,
  output 				       I2C1_SDA_O,
  output 				       I2C1_SDA_T,
  input 				       I2C1_SCL_I,
  output 				       I2C1_SCL_O,
  output 				       I2C1_SCL_T,
  
  //FMIO PJTAG
  input 				       PJTAG_TCK,
  input 				       PJTAG_TMS,
  input 				       PJTAG_TDI,
  output 				       PJTAG_TDO,

  
  //FMIO SDIO0
  output 				       SDIO0_CLK,
  input 				       SDIO0_CLK_FB,
  output 				       SDIO0_CMD_O,
  input 				       SDIO0_CMD_I,
  output 				       SDIO0_CMD_T,
  input [3:0] 				       SDIO0_DATA_I,
  output [3:0] 				       SDIO0_DATA_O,
  output [3:0] 				       SDIO0_DATA_T,
  output 				       SDIO0_LED,
  input 				       SDIO0_CDN,
  input 				       SDIO0_WP, 
  output 				       SDIO0_BUSPOW,
  output [2:0] 				       SDIO0_BUSVOLT,

  //FMIO SDIO1
  output 				       SDIO1_CLK,
  input 				       SDIO1_CLK_FB,
  output 				       SDIO1_CMD_O,
  input 				       SDIO1_CMD_I,
  output 				       SDIO1_CMD_T,
  input [3:0] 				       SDIO1_DATA_I,
  output [3:0] 				       SDIO1_DATA_O,
  output [3:0] 				       SDIO1_DATA_T, 
  output 				       SDIO1_LED,
  input 				       SDIO1_CDN, 
  input 				       SDIO1_WP,
  output 				       SDIO1_BUSPOW, 
  output [2:0] 				       SDIO1_BUSVOLT,

  //FMIO SPI0
  input 				       SPI0_SCLK_I,
  output 				       SPI0_SCLK_O,
  output 				       SPI0_SCLK_T,
  input 				       SPI0_MOSI_I,
  output 				       SPI0_MOSI_O,
  output 				       SPI0_MOSI_T,
  input 				       SPI0_MISO_I,
  output 				       SPI0_MISO_O,
  output 				       SPI0_MISO_T,
  input 				       SPI0_SS_I,
  output 				       SPI0_SS_O,
  output 				       SPI0_SS1_O,
  output 				       SPI0_SS2_O,
  output 				       SPI0_SS_T,

  //FMIO SPI1
  input 				       SPI1_SCLK_I,
  output 				       SPI1_SCLK_O,
  output 				       SPI1_SCLK_T,
  input 				       SPI1_MOSI_I,
  output 				       SPI1_MOSI_O,
  output 				       SPI1_MOSI_T,
  input 				       SPI1_MISO_I,
  output 				       SPI1_MISO_O,
  output 				       SPI1_MISO_T,
  input 				       SPI1_SS_I,
  output 				       SPI1_SS_O,
  output 				       SPI1_SS1_O,
  output 				       SPI1_SS2_O, 
  output 				       SPI1_SS_T,

  //FMIO UART0
  output 				       UART0_DTRN,
  output 				       UART0_RTSN, 
  output 				       UART0_TX,
  input 				       UART0_CTSN,
  input 				       UART0_DCDN,
  input 				       UART0_DSRN,
  input 				       UART0_RIN, 
  input 				       UART0_RX,

  //FMIO UART1
  output 				       UART1_DTRN,
  output 				       UART1_RTSN, 
  output 				       UART1_TX,
  input 				       UART1_CTSN,
  input 				       UART1_DCDN,
  input 				       UART1_DSRN,
  input 				       UART1_RIN, 
  input 				       UART1_RX,

  //FMIO TTC0
  output 				       TTC0_WAVE0_OUT,
  output 				       TTC0_WAVE1_OUT,
  output 				       TTC0_WAVE2_OUT,
  input 				       TTC0_CLK0_IN,
  input 				       TTC0_CLK1_IN,
  input 				       TTC0_CLK2_IN,

  //FMIO TTC1
  output 				       TTC1_WAVE0_OUT,
  output 				       TTC1_WAVE1_OUT,
  output 				       TTC1_WAVE2_OUT,
  input 				       TTC1_CLK0_IN,
  input 				       TTC1_CLK1_IN,
  input 				       TTC1_CLK2_IN,

  //WDT
  input 				       WDT_CLK_IN,
  output 				       WDT_RST_OUT,

  //FTPORT
  input 				       TRACE_CLK,
  output 				       TRACE_CTL,
  output [(C_TRACE_INTERNAL_WIDTH)-1:0]        TRACE_DATA,
  output reg 				       TRACE_CLK_OUT,
  
  // USB
  output [1:0] 				       USB0_PORT_INDCTL,
  output 				       USB0_VBUS_PWRSELECT,
  input 				       USB0_VBUS_PWRFAULT,

  output [1:0] 				       USB1_PORT_INDCTL,
  output 				       USB1_VBUS_PWRSELECT,
  input 				       USB1_VBUS_PWRFAULT,
  
  input 				       SRAM_INTIN,

  //AIO ===================================================

  //M_AXI_GP0
  
  // -- Output
  
  output 				       M_AXI_GP0_ARESETN,
  output 				       M_AXI_GP0_ARVALID,
  output 				       M_AXI_GP0_AWVALID,
  output 				       M_AXI_GP0_BREADY,
  output 				       M_AXI_GP0_RREADY,
  output 				       M_AXI_GP0_WLAST,
  output 				       M_AXI_GP0_WVALID,
  output [(C_M_AXI_GP0_THREAD_ID_WIDTH - 1):0] M_AXI_GP0_ARID,
  output [(C_M_AXI_GP0_THREAD_ID_WIDTH - 1):0] M_AXI_GP0_AWID,
  output [(C_M_AXI_GP0_THREAD_ID_WIDTH - 1):0] M_AXI_GP0_WID,
  output [1:0] 				       M_AXI_GP0_ARBURST,
  output [1:0] 				       M_AXI_GP0_ARLOCK,
  output [2:0] 				       M_AXI_GP0_ARSIZE,
  output [1:0] 				       M_AXI_GP0_AWBURST,
  output [1:0] 				       M_AXI_GP0_AWLOCK,
  output [2:0] 				       M_AXI_GP0_AWSIZE,
  output [2:0] 				       M_AXI_GP0_ARPROT,
  output [2:0] 				       M_AXI_GP0_AWPROT,
  output [31:0] 			       M_AXI_GP0_ARADDR,
  output [31:0] 			       M_AXI_GP0_AWADDR,
  output [31:0] 			       M_AXI_GP0_WDATA,
  output [3:0] 				       M_AXI_GP0_ARCACHE,
  output [3:0] 				       M_AXI_GP0_ARLEN,
  output [3:0] 				       M_AXI_GP0_ARQOS,
  output [3:0] 				       M_AXI_GP0_AWCACHE,
  output [3:0] 				       M_AXI_GP0_AWLEN,
  output [3:0] 				       M_AXI_GP0_AWQOS,
  output [3:0] 				       M_AXI_GP0_WSTRB, 
  
  // -- Input  
  
  input 				       M_AXI_GP0_ACLK,
  input 				       M_AXI_GP0_ARREADY,
  input 				       M_AXI_GP0_AWREADY,
  input 				       M_AXI_GP0_BVALID,
  input 				       M_AXI_GP0_RLAST,
  input 				       M_AXI_GP0_RVALID,
  input 				       M_AXI_GP0_WREADY,
  input [(C_M_AXI_GP0_THREAD_ID_WIDTH - 1):0]  M_AXI_GP0_BID,
  input [(C_M_AXI_GP0_THREAD_ID_WIDTH - 1):0]  M_AXI_GP0_RID,
  input [1:0] 				       M_AXI_GP0_BRESP,
  input [1:0] 				       M_AXI_GP0_RRESP,
  input [31:0] 				       M_AXI_GP0_RDATA, 


  //M_AXI_GP1
  
  // -- Output

  output 				       M_AXI_GP1_ARESETN,
  output 				       M_AXI_GP1_ARVALID,
  output 				       M_AXI_GP1_AWVALID,
  output 				       M_AXI_GP1_BREADY,
  output 				       M_AXI_GP1_RREADY,
  output 				       M_AXI_GP1_WLAST,
  output 				       M_AXI_GP1_WVALID,
  output [(C_M_AXI_GP1_THREAD_ID_WIDTH - 1):0] M_AXI_GP1_ARID,
  output [(C_M_AXI_GP1_THREAD_ID_WIDTH - 1):0] M_AXI_GP1_AWID,
  output [(C_M_AXI_GP1_THREAD_ID_WIDTH - 1):0] M_AXI_GP1_WID,
  output [1:0] 				       M_AXI_GP1_ARBURST,
  output [1:0] 				       M_AXI_GP1_ARLOCK,
  output [2:0] 				       M_AXI_GP1_ARSIZE,
  output [1:0] 				       M_AXI_GP1_AWBURST,
  output [1:0] 				       M_AXI_GP1_AWLOCK,
  output [2:0] 				       M_AXI_GP1_AWSIZE,
  output [2:0] 				       M_AXI_GP1_ARPROT,
  output [2:0] 				       M_AXI_GP1_AWPROT,
  output [31:0] 			       M_AXI_GP1_ARADDR,
  output [31:0] 			       M_AXI_GP1_AWADDR,
  output [31:0] 			       M_AXI_GP1_WDATA,
  output [3:0] 				       M_AXI_GP1_ARCACHE,
  output [3:0] 				       M_AXI_GP1_ARLEN,
  output [3:0] 				       M_AXI_GP1_ARQOS,
  output [3:0] 				       M_AXI_GP1_AWCACHE,
  output [3:0] 				       M_AXI_GP1_AWLEN,
  output [3:0] 				       M_AXI_GP1_AWQOS,
  output [3:0] 				       M_AXI_GP1_WSTRB,
  
  // -- Input
  
  input 				       M_AXI_GP1_ACLK,
  input 				       M_AXI_GP1_ARREADY,
  input 				       M_AXI_GP1_AWREADY,
  input 				       M_AXI_GP1_BVALID,
  input 				       M_AXI_GP1_RLAST,
  input 				       M_AXI_GP1_RVALID,
  input 				       M_AXI_GP1_WREADY, 
  input [(C_M_AXI_GP1_THREAD_ID_WIDTH - 1):0]  M_AXI_GP1_BID,
  input [(C_M_AXI_GP1_THREAD_ID_WIDTH - 1):0]  M_AXI_GP1_RID,
  input [1:0] 				       M_AXI_GP1_BRESP,
  input [1:0] 				       M_AXI_GP1_RRESP,
  input [31:0] 				       M_AXI_GP1_RDATA, 
  

  // S_AXI_GP0
  
  // -- Output
  
  output 				       S_AXI_GP0_ARESETN,
  output 				       S_AXI_GP0_ARREADY,
  output 				       S_AXI_GP0_AWREADY,
  output 				       S_AXI_GP0_BVALID,
  output 				       S_AXI_GP0_RLAST,
  output 				       S_AXI_GP0_RVALID,
  output 				       S_AXI_GP0_WREADY, 
  output [1:0] 				       S_AXI_GP0_BRESP,
  output [1:0] 				       S_AXI_GP0_RRESP,
  output [31:0] 			       S_AXI_GP0_RDATA,
  output [(C_S_AXI_GP0_ID_WIDTH - 1) : 0]      S_AXI_GP0_BID,
  output [(C_S_AXI_GP0_ID_WIDTH - 1) : 0]      S_AXI_GP0_RID,
  
  // -- Input
  input 				       S_AXI_GP0_ACLK,
  input 				       S_AXI_GP0_ARVALID,
  input 				       S_AXI_GP0_AWVALID,
  input 				       S_AXI_GP0_BREADY,
  input 				       S_AXI_GP0_RREADY,
  input 				       S_AXI_GP0_WLAST,
  input 				       S_AXI_GP0_WVALID,
  input [1:0] 				       S_AXI_GP0_ARBURST,
  input [1:0] 				       S_AXI_GP0_ARLOCK,
  input [2:0] 				       S_AXI_GP0_ARSIZE,
  input [1:0] 				       S_AXI_GP0_AWBURST,
  input [1:0] 				       S_AXI_GP0_AWLOCK,
  input [2:0] 				       S_AXI_GP0_AWSIZE,
  input [2:0] 				       S_AXI_GP0_ARPROT,
  input [2:0] 				       S_AXI_GP0_AWPROT,
  input [31:0] 				       S_AXI_GP0_ARADDR,
  input [31:0] 				       S_AXI_GP0_AWADDR,
  input [31:0] 				       S_AXI_GP0_WDATA,
  input [3:0] 				       S_AXI_GP0_ARCACHE,
  input [3:0] 				       S_AXI_GP0_ARLEN,
  input [3:0] 				       S_AXI_GP0_ARQOS,
  input [3:0] 				       S_AXI_GP0_AWCACHE,
  input [3:0] 				       S_AXI_GP0_AWLEN,
  input [3:0] 				       S_AXI_GP0_AWQOS,
  input [3:0] 				       S_AXI_GP0_WSTRB,
  input [(C_S_AXI_GP0_ID_WIDTH - 1) : 0]       S_AXI_GP0_ARID,
  input [(C_S_AXI_GP0_ID_WIDTH - 1) : 0]       S_AXI_GP0_AWID,
  input [(C_S_AXI_GP0_ID_WIDTH - 1) : 0]       S_AXI_GP0_WID, 

  // S_AXI_GP1
  
  // -- Output  
  output 				       S_AXI_GP1_ARESETN,
  output 				       S_AXI_GP1_ARREADY,
  output 				       S_AXI_GP1_AWREADY,
  output 				       S_AXI_GP1_BVALID,
  output 				       S_AXI_GP1_RLAST,
  output 				       S_AXI_GP1_RVALID,
  output 				       S_AXI_GP1_WREADY, 
  output [1:0] 				       S_AXI_GP1_BRESP,
  output [1:0] 				       S_AXI_GP1_RRESP,
  output [31:0] 			       S_AXI_GP1_RDATA,
  output [(C_S_AXI_GP1_ID_WIDTH - 1) : 0]      S_AXI_GP1_BID,
  output [(C_S_AXI_GP1_ID_WIDTH - 1) : 0]      S_AXI_GP1_RID,
  
  // -- Input
  input 				       S_AXI_GP1_ACLK,
  input 				       S_AXI_GP1_ARVALID,
  input 				       S_AXI_GP1_AWVALID,
  input 				       S_AXI_GP1_BREADY,
  input 				       S_AXI_GP1_RREADY,
  input 				       S_AXI_GP1_WLAST,
  input 				       S_AXI_GP1_WVALID,
  input [1:0] 				       S_AXI_GP1_ARBURST,
  input [1:0] 				       S_AXI_GP1_ARLOCK,
  input [2:0] 				       S_AXI_GP1_ARSIZE,
  input [1:0] 				       S_AXI_GP1_AWBURST,
  input [1:0] 				       S_AXI_GP1_AWLOCK,
  input [2:0] 				       S_AXI_GP1_AWSIZE,
  input [2:0] 				       S_AXI_GP1_ARPROT,
  input [2:0] 				       S_AXI_GP1_AWPROT,
  input [31:0] 				       S_AXI_GP1_ARADDR,
  input [31:0] 				       S_AXI_GP1_AWADDR,
  input [31:0] 				       S_AXI_GP1_WDATA,
  input [3:0] 				       S_AXI_GP1_ARCACHE,
  input [3:0] 				       S_AXI_GP1_ARLEN,
  input [3:0] 				       S_AXI_GP1_ARQOS,
  input [3:0] 				       S_AXI_GP1_AWCACHE,
  input [3:0] 				       S_AXI_GP1_AWLEN,
  input [3:0] 				       S_AXI_GP1_AWQOS,
  input [3:0] 				       S_AXI_GP1_WSTRB,
  input [(C_S_AXI_GP1_ID_WIDTH - 1) : 0]       S_AXI_GP1_ARID,
  input [(C_S_AXI_GP1_ID_WIDTH - 1) : 0]       S_AXI_GP1_AWID,
  input [(C_S_AXI_GP1_ID_WIDTH - 1) : 0]       S_AXI_GP1_WID, 

  //S_AXI_ACP
  
  // -- Output  
  
  output 				       S_AXI_ACP_ARESETN,
  output 				       S_AXI_ACP_ARREADY,
  output 				       S_AXI_ACP_AWREADY,
  output 				       S_AXI_ACP_BVALID,
  output 				       S_AXI_ACP_RLAST,
  output 				       S_AXI_ACP_RVALID,
  output 				       S_AXI_ACP_WREADY, 
  output [1:0] 				       S_AXI_ACP_BRESP,
  output [1:0] 				       S_AXI_ACP_RRESP,
  output [(C_S_AXI_ACP_ID_WIDTH - 1) : 0]      S_AXI_ACP_BID,
  output [(C_S_AXI_ACP_ID_WIDTH - 1) : 0]      S_AXI_ACP_RID,
  output [63:0] 			       S_AXI_ACP_RDATA,
  
  // -- Input
  
  input 				       S_AXI_ACP_ACLK,
  input 				       S_AXI_ACP_ARVALID,
  input 				       S_AXI_ACP_AWVALID,
  input 				       S_AXI_ACP_BREADY,
  input 				       S_AXI_ACP_RREADY,
  input 				       S_AXI_ACP_WLAST,
  input 				       S_AXI_ACP_WVALID,
  input [(C_S_AXI_ACP_ID_WIDTH - 1) : 0]       S_AXI_ACP_ARID,
  input [2:0] 				       S_AXI_ACP_ARPROT,
  input [(C_S_AXI_ACP_ID_WIDTH - 1) : 0]       S_AXI_ACP_AWID,
  input [2:0] 				       S_AXI_ACP_AWPROT,
  input [(C_S_AXI_ACP_ID_WIDTH - 1) : 0]       S_AXI_ACP_WID,
  input [31:0] 				       S_AXI_ACP_ARADDR,
  input [31:0] 				       S_AXI_ACP_AWADDR,
  input [3:0] 				       S_AXI_ACP_ARCACHE,
  input [3:0] 				       S_AXI_ACP_ARLEN,
  input [3:0] 				       S_AXI_ACP_ARQOS,
  input [3:0] 				       S_AXI_ACP_AWCACHE,
  input [3:0] 				       S_AXI_ACP_AWLEN,
  input [3:0] 				       S_AXI_ACP_AWQOS, 
  input [1:0] 				       S_AXI_ACP_ARBURST,
  input [1:0] 				       S_AXI_ACP_ARLOCK,
  input [2:0] 				       S_AXI_ACP_ARSIZE,
  input [1:0] 				       S_AXI_ACP_AWBURST,
  input [1:0] 				       S_AXI_ACP_AWLOCK,
  input [2:0] 				       S_AXI_ACP_AWSIZE,
  input [4:0] 				       S_AXI_ACP_ARUSER,
  input [4:0] 				       S_AXI_ACP_AWUSER,
  input [63:0] 				       S_AXI_ACP_WDATA,
  input [7:0] 				       S_AXI_ACP_WSTRB, 
  
  // S_AXI_HP_0
  
  // -- Output
  output 				       S_AXI_HP0_ARESETN,
  output 				       S_AXI_HP0_ARREADY,
  output 				       S_AXI_HP0_AWREADY,
  output 				       S_AXI_HP0_BVALID,
  output 				       S_AXI_HP0_RLAST,
  output 				       S_AXI_HP0_RVALID,
  output 				       S_AXI_HP0_WREADY, 
  output [1:0] 				       S_AXI_HP0_BRESP,
  output [1:0] 				       S_AXI_HP0_RRESP,
  output [(C_S_AXI_HP0_ID_WIDTH - 1) : 0]      S_AXI_HP0_BID,
  output [(C_S_AXI_HP0_ID_WIDTH - 1) : 0]      S_AXI_HP0_RID,
  output [(C_S_AXI_HP0_DATA_WIDTH - 1) :0]     S_AXI_HP0_RDATA,
  output [7:0] 				       S_AXI_HP0_RCOUNT,
  output [7:0] 				       S_AXI_HP0_WCOUNT,
  output [2:0] 				       S_AXI_HP0_RACOUNT,
  output [5:0] 				       S_AXI_HP0_WACOUNT,
  
  // -- Input  
  input 				       S_AXI_HP0_ACLK,
  input 				       S_AXI_HP0_ARVALID,
  input 				       S_AXI_HP0_AWVALID,
  input 				       S_AXI_HP0_BREADY,
  input 				       S_AXI_HP0_RDISSUECAP1_EN,
  input 				       S_AXI_HP0_RREADY,
  input 				       S_AXI_HP0_WLAST,
  input 				       S_AXI_HP0_WRISSUECAP1_EN,
  input 				       S_AXI_HP0_WVALID,
  input [1:0] 				       S_AXI_HP0_ARBURST,
  input [1:0] 				       S_AXI_HP0_ARLOCK,
  input [2:0] 				       S_AXI_HP0_ARSIZE,
  input [1:0] 				       S_AXI_HP0_AWBURST,
  input [1:0] 				       S_AXI_HP0_AWLOCK,
  input [2:0] 				       S_AXI_HP0_AWSIZE,
  input [2:0] 				       S_AXI_HP0_ARPROT,
  input [2:0] 				       S_AXI_HP0_AWPROT,
  input [31:0] 				       S_AXI_HP0_ARADDR,
  input [31:0] 				       S_AXI_HP0_AWADDR,
  input [3:0] 				       S_AXI_HP0_ARCACHE,
  input [3:0] 				       S_AXI_HP0_ARLEN,
  input [3:0] 				       S_AXI_HP0_ARQOS,
  input [3:0] 				       S_AXI_HP0_AWCACHE,
  input [3:0] 				       S_AXI_HP0_AWLEN,
  input [3:0] 				       S_AXI_HP0_AWQOS,
  input [(C_S_AXI_HP0_ID_WIDTH - 1) : 0]       S_AXI_HP0_ARID,
  input [(C_S_AXI_HP0_ID_WIDTH - 1) : 0]       S_AXI_HP0_AWID,
  input [(C_S_AXI_HP0_ID_WIDTH - 1) : 0]       S_AXI_HP0_WID,
  input [(C_S_AXI_HP0_DATA_WIDTH - 1) :0]      S_AXI_HP0_WDATA,
  input [((C_S_AXI_HP0_DATA_WIDTH/8)-1):0]     S_AXI_HP0_WSTRB, 

  // S_AXI_HP1
  // -- Output
  output 				       S_AXI_HP1_ARESETN,
  output 				       S_AXI_HP1_ARREADY,
  output 				       S_AXI_HP1_AWREADY,
  output 				       S_AXI_HP1_BVALID,
  output 				       S_AXI_HP1_RLAST,
  output 				       S_AXI_HP1_RVALID,
  output 				       S_AXI_HP1_WREADY, 
  output [1:0] 				       S_AXI_HP1_BRESP,
  output [1:0] 				       S_AXI_HP1_RRESP,
  output [(C_S_AXI_HP1_ID_WIDTH - 1) : 0]      S_AXI_HP1_BID,
  output [(C_S_AXI_HP1_ID_WIDTH - 1) : 0]      S_AXI_HP1_RID,
  output [(C_S_AXI_HP1_DATA_WIDTH - 1) :0]     S_AXI_HP1_RDATA,
  output [7:0] 				       S_AXI_HP1_RCOUNT,
  output [7:0] 				       S_AXI_HP1_WCOUNT,
  output [2:0] 				       S_AXI_HP1_RACOUNT,
  output [5:0] 				       S_AXI_HP1_WACOUNT,
  
  
  // -- Input  
  input 				       S_AXI_HP1_ACLK,
  input 				       S_AXI_HP1_ARVALID,
  input 				       S_AXI_HP1_AWVALID,
  input 				       S_AXI_HP1_BREADY,
  input 				       S_AXI_HP1_RDISSUECAP1_EN,
  input 				       S_AXI_HP1_RREADY,
  input 				       S_AXI_HP1_WLAST,
  input 				       S_AXI_HP1_WRISSUECAP1_EN,
  input 				       S_AXI_HP1_WVALID,
  input [1:0] 				       S_AXI_HP1_ARBURST,
  input [1:0] 				       S_AXI_HP1_ARLOCK,
  input [2:0] 				       S_AXI_HP1_ARSIZE,
  input [1:0] 				       S_AXI_HP1_AWBURST,
  input [1:0] 				       S_AXI_HP1_AWLOCK,
  input [2:0] 				       S_AXI_HP1_AWSIZE,
  input [2:0] 				       S_AXI_HP1_ARPROT,
  input [2:0] 				       S_AXI_HP1_AWPROT,
  input [31:0] 				       S_AXI_HP1_ARADDR,
  input [31:0] 				       S_AXI_HP1_AWADDR,
  input [3:0] 				       S_AXI_HP1_ARCACHE,
  input [3:0] 				       S_AXI_HP1_ARLEN,
  input [3:0] 				       S_AXI_HP1_ARQOS,
  input [3:0] 				       S_AXI_HP1_AWCACHE,
  input [3:0] 				       S_AXI_HP1_AWLEN,
  input [3:0] 				       S_AXI_HP1_AWQOS,
  input [(C_S_AXI_HP1_ID_WIDTH - 1) : 0]       S_AXI_HP1_ARID,
  input [(C_S_AXI_HP1_ID_WIDTH - 1) : 0]       S_AXI_HP1_AWID,
  input [(C_S_AXI_HP1_ID_WIDTH - 1) : 0]       S_AXI_HP1_WID,
  input [(C_S_AXI_HP1_DATA_WIDTH - 1) :0]      S_AXI_HP1_WDATA,
  input [((C_S_AXI_HP1_DATA_WIDTH/8)-1):0]     S_AXI_HP1_WSTRB, 

  // S_AXI_HP2
  // -- Output
  output 				       S_AXI_HP2_ARESETN,
  output 				       S_AXI_HP2_ARREADY,
  output 				       S_AXI_HP2_AWREADY,
  output 				       S_AXI_HP2_BVALID,
  output 				       S_AXI_HP2_RLAST,
  output 				       S_AXI_HP2_RVALID,
  output 				       S_AXI_HP2_WREADY, 
  output [1:0] 				       S_AXI_HP2_BRESP,
  output [1:0] 				       S_AXI_HP2_RRESP,
  output [(C_S_AXI_HP2_ID_WIDTH - 1) : 0]      S_AXI_HP2_BID,
  output [(C_S_AXI_HP2_ID_WIDTH - 1) : 0]      S_AXI_HP2_RID,
  output [(C_S_AXI_HP2_DATA_WIDTH - 1) :0]     S_AXI_HP2_RDATA,
  output [7:0] 				       S_AXI_HP2_RCOUNT,
  output [7:0] 				       S_AXI_HP2_WCOUNT,
  output [2:0] 				       S_AXI_HP2_RACOUNT,
  output [5:0] 				       S_AXI_HP2_WACOUNT,
  
  
  // -- Input  
  input 				       S_AXI_HP2_ACLK,
  input 				       S_AXI_HP2_ARVALID,
  input 				       S_AXI_HP2_AWVALID,
  input 				       S_AXI_HP2_BREADY,
  input 				       S_AXI_HP2_RDISSUECAP1_EN,
  input 				       S_AXI_HP2_RREADY,
  input 				       S_AXI_HP2_WLAST,
  input 				       S_AXI_HP2_WRISSUECAP1_EN,
  input 				       S_AXI_HP2_WVALID,
  input [1:0] 				       S_AXI_HP2_ARBURST,
  input [1:0] 				       S_AXI_HP2_ARLOCK,
  input [2:0] 				       S_AXI_HP2_ARSIZE,
  input [1:0] 				       S_AXI_HP2_AWBURST,
  input [1:0] 				       S_AXI_HP2_AWLOCK,
  input [2:0] 				       S_AXI_HP2_AWSIZE,
  input [2:0] 				       S_AXI_HP2_ARPROT,
  input [2:0] 				       S_AXI_HP2_AWPROT,
  input [31:0] 				       S_AXI_HP2_ARADDR,
  input [31:0] 				       S_AXI_HP2_AWADDR,
  input [3:0] 				       S_AXI_HP2_ARCACHE,
  input [3:0] 				       S_AXI_HP2_ARLEN,
  input [3:0] 				       S_AXI_HP2_ARQOS,
  input [3:0] 				       S_AXI_HP2_AWCACHE,
  input [3:0] 				       S_AXI_HP2_AWLEN,
  input [3:0] 				       S_AXI_HP2_AWQOS,
  input [(C_S_AXI_HP2_ID_WIDTH - 1) : 0]       S_AXI_HP2_ARID,
  input [(C_S_AXI_HP2_ID_WIDTH - 1) : 0]       S_AXI_HP2_AWID,
  input [(C_S_AXI_HP2_ID_WIDTH - 1) : 0]       S_AXI_HP2_WID,
  input [(C_S_AXI_HP2_DATA_WIDTH - 1) :0]      S_AXI_HP2_WDATA,
  input [((C_S_AXI_HP2_DATA_WIDTH/8)-1):0]     S_AXI_HP2_WSTRB, 

  // S_AXI_HP_3
  
  // -- Output
  output 				       S_AXI_HP3_ARESETN,
  output 				       S_AXI_HP3_ARREADY,
  output 				       S_AXI_HP3_AWREADY,
  output 				       S_AXI_HP3_BVALID,
  output 				       S_AXI_HP3_RLAST,
  output 				       S_AXI_HP3_RVALID,
  output 				       S_AXI_HP3_WREADY, 
  output [1:0] 				       S_AXI_HP3_BRESP,
  output [1:0] 				       S_AXI_HP3_RRESP,
  output [(C_S_AXI_HP3_ID_WIDTH - 1) : 0]      S_AXI_HP3_BID,
  output [(C_S_AXI_HP3_ID_WIDTH - 1) : 0]      S_AXI_HP3_RID,
  output [(C_S_AXI_HP3_DATA_WIDTH - 1) :0]     S_AXI_HP3_RDATA,
  output [7:0] 				       S_AXI_HP3_RCOUNT,
  output [7:0] 				       S_AXI_HP3_WCOUNT,
  output [2:0] 				       S_AXI_HP3_RACOUNT,
  output [5:0] 				       S_AXI_HP3_WACOUNT,
  
  
  // -- Input  
  input 				       S_AXI_HP3_ACLK,
  input 				       S_AXI_HP3_ARVALID,
  input 				       S_AXI_HP3_AWVALID,
  input 				       S_AXI_HP3_BREADY,
  input 				       S_AXI_HP3_RDISSUECAP1_EN,
  input 				       S_AXI_HP3_RREADY,
  input 				       S_AXI_HP3_WLAST,
  input 				       S_AXI_HP3_WRISSUECAP1_EN,
  input 				       S_AXI_HP3_WVALID,
  input [1:0] 				       S_AXI_HP3_ARBURST,
  input [1:0] 				       S_AXI_HP3_ARLOCK,
  input [2:0] 				       S_AXI_HP3_ARSIZE,
  input [1:0] 				       S_AXI_HP3_AWBURST,
  input [1:0] 				       S_AXI_HP3_AWLOCK,
  input [2:0] 				       S_AXI_HP3_AWSIZE,
  input [2:0] 				       S_AXI_HP3_ARPROT,
  input [2:0] 				       S_AXI_HP3_AWPROT,
  input [31:0] 				       S_AXI_HP3_ARADDR,
  input [31:0] 				       S_AXI_HP3_AWADDR,
  input [3:0] 				       S_AXI_HP3_ARCACHE,
  input [3:0] 				       S_AXI_HP3_ARLEN,
  input [3:0] 				       S_AXI_HP3_ARQOS,
  input [3:0] 				       S_AXI_HP3_AWCACHE,
  input [3:0] 				       S_AXI_HP3_AWLEN,
  input [3:0] 				       S_AXI_HP3_AWQOS,
  input [(C_S_AXI_HP3_ID_WIDTH - 1) : 0]       S_AXI_HP3_ARID,
  input [(C_S_AXI_HP3_ID_WIDTH - 1) : 0]       S_AXI_HP3_AWID,
  input [(C_S_AXI_HP3_ID_WIDTH - 1) : 0]       S_AXI_HP3_WID,
  input [(C_S_AXI_HP3_DATA_WIDTH - 1) :0]      S_AXI_HP3_WDATA,
  input [((C_S_AXI_HP3_DATA_WIDTH/8)-1):0]     S_AXI_HP3_WSTRB, 
  
  //FIO ========================================

  //IRQ
  output 				       IRQ_P2F_DMAC_ABORT ,
  output 				       IRQ_P2F_DMAC0,
  output 				       IRQ_P2F_DMAC1,
  output 				       IRQ_P2F_DMAC2,
  output 				       IRQ_P2F_DMAC3,
  output 				       IRQ_P2F_DMAC4,
  output 				       IRQ_P2F_DMAC5,
  output 				       IRQ_P2F_DMAC6,
  output 				       IRQ_P2F_DMAC7,
  output 				       IRQ_P2F_SMC,
  output 				       IRQ_P2F_QSPI,
  output 				       IRQ_P2F_CTI,
  output 				       IRQ_P2F_GPIO,
  output 				       IRQ_P2F_USB0,
  output 				       IRQ_P2F_ENET0,
  output 				       IRQ_P2F_ENET_WAKE0,
  output 				       IRQ_P2F_SDIO0,
  output 				       IRQ_P2F_I2C0,
  output 				       IRQ_P2F_SPI0,
  output 				       IRQ_P2F_UART0,
  output 				       IRQ_P2F_CAN0,
  output 				       IRQ_P2F_USB1,
  output 				       IRQ_P2F_ENET1,
  output 				       IRQ_P2F_ENET_WAKE1,
  output 				       IRQ_P2F_SDIO1,
  output 				       IRQ_P2F_I2C1,
  output 				       IRQ_P2F_SPI1,
  output 				       IRQ_P2F_UART1,
  output 				       IRQ_P2F_CAN1,
  input [(C_NUM_F2P_INTR_INPUTS-1):0] 	       IRQ_F2P,
  input 				       Core0_nFIQ,
  input 				       Core0_nIRQ,
  input 				       Core1_nFIQ,
  input 				       Core1_nIRQ,

  //DMA

  output [1:0] 				       DMA0_DATYPE, 
  output 				       DMA0_DAVALID,
  output 				       DMA0_DRREADY,
  output 				       DMA0_RSTN, 
  output [1:0] 				       DMA1_DATYPE, 
  output 				       DMA1_DAVALID,
  output 				       DMA1_DRREADY,
  output 				       DMA1_RSTN, 
  output [1:0] 				       DMA2_DATYPE, 
  output 				       DMA2_DAVALID,
  output 				       DMA2_DRREADY,
  output 				       DMA2_RSTN, 
  output [1:0] 				       DMA3_DATYPE, 
  output 				       DMA3_DAVALID,
  output 				       DMA3_DRREADY,
  output 				       DMA3_RSTN, 
  input 				       DMA0_ACLK,
  input 				       DMA0_DAREADY,
  input 				       DMA0_DRLAST,
  input 				       DMA0_DRVALID,
  input 				       DMA1_ACLK,
  input 				       DMA1_DAREADY,
  input 				       DMA1_DRLAST,
  input 				       DMA1_DRVALID,
  input 				       DMA2_ACLK,
  input 				       DMA2_DAREADY,
  input 				       DMA2_DRLAST,
  input 				       DMA2_DRVALID,
  input 				       DMA3_ACLK,
  input 				       DMA3_DAREADY,
  input 				       DMA3_DRLAST,
  input 				       DMA3_DRVALID, 
  input [1:0] 				       DMA0_DRTYPE,
  input [1:0] 				       DMA1_DRTYPE,
  input [1:0] 				       DMA2_DRTYPE,
  input [1:0] 				       DMA3_DRTYPE,
  
  //FCLK
  output 				       FCLK_CLK3,
  output 				       FCLK_CLK2,
  output 				       FCLK_CLK1,
  output 				       FCLK_CLK0,
 
  input 				       FCLK_CLKTRIG3_N,
  input 				       FCLK_CLKTRIG2_N,
  input 				       FCLK_CLKTRIG1_N,
  input 				       FCLK_CLKTRIG0_N,
 
  output 				       FCLK_RESET3_N,
  output 				       FCLK_RESET2_N,
  output 				       FCLK_RESET1_N,
  output 				       FCLK_RESET0_N,

  //FTMD
  input [31:0] 				       FTMD_TRACEIN_DATA,
  input 				       FTMD_TRACEIN_VALID,
  input 				       FTMD_TRACEIN_CLK,
  input [3:0] 				       FTMD_TRACEIN_ATID,

  //FTMT
  input 				       FTMT_F2P_TRIG_0,
  output 				       FTMT_F2P_TRIGACK_0,
  input 				       FTMT_F2P_TRIG_1,
  output 				       FTMT_F2P_TRIGACK_1,
  input 				       FTMT_F2P_TRIG_2,
  output 				       FTMT_F2P_TRIGACK_2,
  input 				       FTMT_F2P_TRIG_3,
  output 				       FTMT_F2P_TRIGACK_3,
  input [31:0] 				       FTMT_F2P_DEBUG, 
  input 				       FTMT_P2F_TRIGACK_0,
  output 				       FTMT_P2F_TRIG_0,
  input 				       FTMT_P2F_TRIGACK_1,
  output 				       FTMT_P2F_TRIG_1,
  input 				       FTMT_P2F_TRIGACK_2,
  output 				       FTMT_P2F_TRIG_2,
  input 				       FTMT_P2F_TRIGACK_3,
  output 				       FTMT_P2F_TRIG_3,
  output [31:0] 			       FTMT_P2F_DEBUG,

  //FIDLE
  input 				       FPGA_IDLE_N,
  
  //EVENT

  output 				       EVENT_EVENTO,
  output [1:0] 				       EVENT_STANDBYWFE,
  output [1:0] 				       EVENT_STANDBYWFI, 
  input 				       EVENT_EVENTI, 
  

  //DARB
  input [3:0] 				       DDR_ARB,
  inout [C_MIO_PRIMITIVE - 1:0] 	       MIO, 
  
  //DDR
  inout 				       DDR_CAS_n, // CASB
  inout 				       DDR_CKE, // CKE
  inout 				       DDR_Clk_n, // CKN
  inout 				       DDR_Clk, // CKP
  inout 				       DDR_CS_n, // CSB 
  inout 				       DDR_DRSTB, // DDR_DRSTB  
  inout 				       DDR_ODT, // ODT
  inout 				       DDR_RAS_n, // RASB
  inout 				       DDR_WEB,
  inout [2:0] 				       DDR_BankAddr, // BA  
  inout [14:0] 				       DDR_Addr, // A
  
  inout 				       DDR_VRN,
  inout 				       DDR_VRP,
  inout [C_DM_WIDTH - 1:0] 		       DDR_DM, // DM  
  inout [C_DQ_WIDTH - 1:0] 		       DDR_DQ, // DQ
  inout [C_DQS_WIDTH -1:0] 		       DDR_DQS_n, // DQSN
  inout [C_DQS_WIDTH - 1:0] 		       DDR_DQS, // DQSP
  
  inout 				       PS_SRSTB, // SRSTB    
  inout 				       PS_CLK, // CLK
  inout 				       PS_PORB         // PORB 

);

endmodule // processing_system7



