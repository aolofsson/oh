module oh_gray2bin (/*AUTOARG*/
   // Outputs
   out,
   // Inputs
   a
   );

   //###############################################################
   //# Interface
   //###############################################################

   parameter DW = 64;

   input [DW-1:0]  a;         //gray encoded input
   output [DW-1:0] out;       //binary output

   //###############################################################
   //# BODY
   //###############################################################

   
   
   
endmodule // oh_gray2bin



