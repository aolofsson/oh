module oh_ser2par (/*AUTOINST*/);

endmodule // oh_pll
