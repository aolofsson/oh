module oh_ecc_write (/*AUTOARG*/);


endmodule // oh_ecc_write

