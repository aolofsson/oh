//#############################################################################
//# Function: 4 Input Or Gate                                                 #
//# Copyright: OH Project Authors. All rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_or4
   (
    input  a,
    input  b,
    input  c,
    input  d,
    output z
    );

   assign z = a | b | c | d;

endmodule
