module oh_bin2gray (/*AUTOARG*/
   // Outputs
   out,
   // Inputs
   a
   );

   //###############################################################
   //# Interface
   //###############################################################

   parameter DW = 64;

   input [DW-1:0]  a;         //binary input
   output [DW-1:0] out;       //gray-encoded output

   //###############################################################
   //# BODY
   //###############################################################

   
   
   
endmodule // oh_bin2gray


