`define CFG_MIOW   8
`define CFG_MIOPW  104
`define CFG_TARGET "GENERIC"
`define CFG_RANDOM "1"
