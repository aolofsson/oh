module oh_par2ser (/*AUTOINST*/);

endmodule // oh_pll
