module oh_pll (/*AUTOINST*/);

endmodule // oh_pll
