`ifndef EMAILBOX_REGMAP_V_
 `define EMAILBOX_REGMAP_V_

 `ifndef EGROUP_MMR
  `define EGROUP_MMR 4'hf
 `endif

  `define REG_INPUT0 6'h0
  `define REG_INPUT1 6'h1
  `define REG_OUTPUT 6'h2

 `endif


