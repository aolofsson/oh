`ifndef MIO_CONSTANTS_V_
 `define MIO_CONSTANTS_V_

 `define CFG_TARGET "GENERIC"  // default hard macro target
                               // see also "XILINX", "ALTERA", "ASIC"
`endif
