//#############################################################################
//# Function: Tie High Cell                                                   #
//# Copyright: OH Project Authors. ALl rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_tiehi
   (
    output z
    );

   assign z = 1'b1;

endmodule
