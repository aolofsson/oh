//#############################################################################
//# Function: Antenna Diode                                                   #
//# Copyright: OH Project Authors. ALl rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_antenna
   (
    input  vss,
    output z
    );

endmodule
