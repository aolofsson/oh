module BUFIO (/*AUTOARG*/
   // Outputs
   O,
   // Inputs
   I
   );
   input I;
   output O;
   
endmodule // BUFIO

