//#############################################################################
//# Function: Tie Low Cell                                                    #
//# Copyright: OH Project Authors. ALl rights Reserved.                       #
//# License:  MIT (see LICENSE file in OH repository)                         #
//#############################################################################

module asic_tielo #(parameter PROP = "DEFAULT")  (
   output z
   );

   assign z = 1'b0;

endmodule
